library verilog;
use verilog.vl_types.all;
entity ula_of_infinity_vlg_vec_tst is
end ula_of_infinity_vlg_vec_tst;
