library verilog;
use verilog.vl_types.all;
entity machine_calc_vlg_vec_tst is
end machine_calc_vlg_vec_tst;
