library verilog;
use verilog.vl_types.all;
entity mux4_1b_vlg_check_tst is
    port(
        \out\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux4_1b_vlg_check_tst;
