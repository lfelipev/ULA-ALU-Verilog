library verilog;
use verilog.vl_types.all;
entity test_machine_vlg_vec_tst is
end test_machine_vlg_vec_tst;
