library verilog;
use verilog.vl_types.all;
entity machine_of_destiny_vlg_vec_tst is
end machine_of_destiny_vlg_vec_tst;
