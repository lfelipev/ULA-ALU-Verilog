library verilog;
use verilog.vl_types.all;
entity mux4_1b_vlg_vec_tst is
end mux4_1b_vlg_vec_tst;
