library verilog;
use verilog.vl_types.all;
entity final_test_machine_vlg_vec_tst is
end final_test_machine_vlg_vec_tst;
