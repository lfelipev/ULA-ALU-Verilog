library verilog;
use verilog.vl_types.all;
entity mux2_1b_vlg_vec_tst is
end mux2_1b_vlg_vec_tst;
